module InstructionMmem (
    input wire [4:0] address,
    output reg [31:0] inst
);

	//reg [31:0] inst;

	always @(address) begin
		case(address)
			00 : inst = 32'h20020005;
			01 : inst = 32'h20070003;
			02 : inst = 32'h2003000c;
			03 : inst = 32'h00e22025;
			04 : inst = 32'h00642824;
			05 : inst = 32'h00a42820;
			06 : inst = 32'h10a70008;
			07 : inst = 32'h0064302a;
			08 : inst = 32'h10c00001;
			09 : inst = 32'h2005000a;
			10 : inst = 32'h00e2302a;
			11 : inst = 32'h00c53820;
			12 : inst = 32'h00e23822;
			13 : inst = 32'h0800000f;
			14 : inst = 32'h8c070000;
			15 : inst = 32'hac470047;
			16 : inst = 32'h00000000;
			17 : inst = 32'h00000000;
			18 : inst = 32'h00000000;
			19 : inst = 32'h00000000;
			20 : inst = 32'h00000000;
			21 : inst = 32'h00000000;
			22 : inst = 32'h00000000;
			23 : inst = 32'h00000000;
			24 : inst = 32'h00000000;
			25 : inst = 32'h00000000;
			26 : inst = 32'h00000000;
			27 : inst = 32'h00000000;
			28 : inst = 32'h00000000;
			29 : inst = 32'h00000000;
			30 : inst = 32'h00000000;
			31 : inst = 32'h00000000;
			32 : inst = 32'h00000000;
			33 : inst = 32'h00000000;
			34 : inst = 32'h00000000;
			35 : inst = 32'h00000000;
			36 : inst = 32'h00000000;
			37 : inst = 32'h00000000;
			38 : inst = 32'h00000000;
			39 : inst = 32'h00000000;
			40 : inst = 32'h00000000;
			41 : inst = 32'h00000000;
			42 : inst = 32'h00000000;
			43 : inst = 32'h00000000;
			44 : inst = 32'h00000000;
			45 : inst = 32'h00000000;
			46 : inst = 32'h00000000;
			47 : inst = 32'h00000000;
			48 : inst = 32'h00000000;
			49 : inst = 32'h00000000;
			50 : inst = 32'h00000000;
			51 : inst = 32'h00000000;
			52 : inst = 32'h00000000;
			53 : inst = 32'h00000000;
			54 : inst = 32'h00000000;
			55 : inst = 32'h00000000;
			56 : inst = 32'h00000000;
			57 : inst = 32'h00000000;
			58 : inst = 32'h00000000;
			59 : inst = 32'h00000000;
			60 : inst = 32'h00000000;
			61 : inst = 32'h00000000;
			62 : inst = 32'h00000000;
			63 : inst = 32'h00000000;
		endcase
	end

endmodule
